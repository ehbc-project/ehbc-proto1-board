library ieee;
use ieee.std_logic_1164.all;

package common is
    -- MEMC/CASGEN/RASGEN Common Type
    type strobe_mode_t is ( SEM_NONE, SEM_SEL, SEM_ALL );
end common;

package body common is
end common;
